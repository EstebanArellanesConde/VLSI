-- PROGRAMA ESTANDAR PARA CARTA FMS Y ASM
-- M.I. BRYAN EMMANUEL ALVAREZ SERNA

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY fsm IS
	PORT(ENTRADAS, CLK: IN STD_LOGIC;
	       SALIDA: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE BEAS OF fsm IS
TYPE ESTADOS IS (INICIO, ESTADO1, ESTADO2);
SIGNAL PRESENTE: ESTADOS := INICIO;
BEGIN

	PROCESS(ENTRADAS,CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			CASE PRESENTE IS
				WHEN INICIO => -- TAREAS EN INICIO
				
				WHEN ESTADO1 => -- TAREAS EN ESTADO1
				
				WHEN ESTADO2 => -- TAREAS EN ESTADO2
				--SE PUEDEN AGREGAR TODOS LOS ESTADOS QUE SE NECESITEN
			END CASE;
		END IF;
	END PROCESS;

END BEAS;
