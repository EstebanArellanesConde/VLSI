LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ffd2 IS 
	PORT ( BOT: IN STD_LOGIC;
		    CLK: IN STD_LOGIC;
			 Q1: BUFFER STD_LOGIC;
		    Q2: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE BEAS OF ffd2 IS
BEGIN

	PROCESS(CLK)
	BEGIN
		IF RISING_EDGE (CLK) THEN 
			Q1 <= BOT;
			Q2 <= Q1;
		END IF;
	END PROCESS;

	
END BEAS;
