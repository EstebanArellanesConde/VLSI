
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY Comp IS
PORT (CT, CUENTA: IN INTEGER RANGE 0 TO 9; CLK: IN STD_LOGIC;
END ENTITY;
PWM: OUT STD_LOGIC);
ARCHITECTURE BEAS OF comp IS
SIGNAL PWMQ: STD_LOGIC;
BEGIN
PROCESS (CUENTA)
BEGIN
IF CUENTA <- CT THEN
PWMQ<= '1';
ELSE
PWMQ <= '0';
END IF;
END PROCESS;
PROCESS (CLK)
BEGIN
IF FALLING EDGE (CLK) THEN
PWM <= PWMQ;
END IF;
END PROCESS;
END BEAS;