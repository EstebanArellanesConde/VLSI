LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX IS
PORT(CLK: IN STD_LOGIC
;
UN, DEC: IN STD_LOGIC_VECTOR (6 downto 0);
D1,D2: OUT STD_LOGIC;
DIG: OUT STD_LOGIC_VECTOR (6 downto 0));

END ENTITY;
ARCHITECTURE ALGO OF MUX IS
SIGNAL AUX2: STD_LOGIC
;

BEGIN

PROCESS(CLK)
BEGIN
IF RISING_EDGE(CLK) THE
N
IF AUX2='1' THEN
D1<='1';
D2<='0';
DIG<=UN;
AUX2<=NOT AUX2;

ELSE

D2<='1';
D1<='0';
DIG<=DEC;
AUX2<=NOT AUX2;

END IF;

END IF;
END PROCESS;
END ALGO;
