LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY conta IS 
	PORT ( RST, CLK: IN STD_LOGIC;)
	
END ENTITY;

ARCHITECTURE BEAS OF conta IS
BEGIN

	PROCESS(CLK)
	BEGIN
		IF RISING_EDGE (CLK) THEN 
			IF CUENTA = '1' THEN
				CUENTA <= 0;
			ELSIF CUENTA = 3 THEN
				CUENTA <= 0;
			ELSE
				CUENTA <= CUENTA + 1;
		END IF;
	END PROCESS;

	
END BEAS;
