LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY contac IS 
	PORT (RST, CLK: IN STD_LOGIC;
		    CARRY: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE ALGO OF contac IS
SIGNAL CUENTA:INTEGER RANGE 0 TO 524287;

BEGIN

			PROCESS (CLK,RST)
			BEGIN 
				IF RST='1' THEN
					CUENTA<=0;
					CARRY<='0';
				ELSIF RISING_EDGE (CLK) THEN
					IF CUENTA=524287 THEN
						CARRY<='1'; 
					ELSE
						CUENTA<=CUENTA+1;
						CARRY<='0';
					END IF;
					
				END IF;
			END PROCESS;

			
END ALGO;
