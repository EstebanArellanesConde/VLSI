-- PROGRAMA ESTANDAR PARA CARTA FMS Y ASM
-- M.I. BRYAN EMMANUEL ALVAREZ SERNA

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY fsm IS
	PORT(BOT, CLK: IN STD_LOGIC;
	       SALIDA: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE BEAS OF fsm IS
TYPE ESTADOS IS (INICIO, ESTADO1, ESTADO2, ESTADO3);
SIGNAL PRESENTE: ESTADOS := INICIO;
BEGIN

	PROCESS(BOT,CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			CASE PRESENTE IS
				WHEN INICIO => -- TAREAS EN INICIO
					SALIDA <= '0';
					IF BOT = '0' THEN
						PRESENTE <= INICIO;
					ELSE
                  PRESENTE <= ESTADO1; -- Cambia a ESTADO1
               END IF;
				WHEN ESTADO1 => -- TAREAS EN ESTADO1
					SALIDA <= '1';
					IF BOT = '1' THEN
						PRESENTE <= ESTADO1;
					ELSE
                  PRESENTE <= ESTADO2;
					END IF;
				WHEN ESTADO2 => -- TAREAS EN ESTADO2
					SALIDA <= '1';
					IF BOT = '0' THEN
						PRESENTE <= ESTADO2;
					ELSE
                  PRESENTE <= ESTADO3;
					END IF;
				WHEN ESTADO3 => -- TAREAS EN ESTADO3
					SALIDA <= '0';
					IF BOT = '1' THEN
						PRESENTE <= ESTADO3;
					ELSE
                  PRESENTE <= INICIO;
					END IF;
				--SE PUEDEN AGREGAR TODOS LOS ESTADOS QUE SE NECESITEN
			END CASE;
		END IF;
	END PROCESS;

END BEAS;
