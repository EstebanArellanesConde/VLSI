LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY CONT99 IS

PORT(CLK, UD, RST: IN STD_LOGIC;
ONE: OUT STD_LOGIC;
CUENTAU,CUENTAD: OUT STD_LOGIC_VECTOR (3 downto 0));

END ENTITY;
ARCHITECTURE ALGO OF CONT99 IS

SIGNAL AUXU,AUXD: STD_LOGIC_VECTOR (3 downto 0);
BEGIN

PROCESS(CLK, RST,UD)
BEGIN

IF (RST='0') THEN

AUXU<="0000";
AUXD<="0000";
ELSIF FALLING_EDGE (CLK) THEN
IF (UD='1') THEN

IF AUXU="1001" THEN
AUXU<= "0000";

IF AUXD="1001" THEN
AUXD<="0000";
ELSE
AUXD<=AUXD+'1';
END IF;

ELSE
AUXU<=AUXU+'1';
END IF;

ELSE

IF AUXU="0000" THEN
AUXU<="1001";

IF AUXD="0000" THEN
AUXD<="1001";
ELSE
AUXD<=AUXD­'1';
END IF;

ELSE
AUXU<=AUXU­'1';
END IF;

END IF;

END IF;
END PROCESS;
CUENTAU<= AUXU;
CUENTAD<=AUXD;
ONE<='1';
END ARCHITECTURE;
