LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ffdh IS 
	PORT ( HAB: IN STD_LOGIC;
	       D: IN STD_LOGIC;
		    CLK: IN STD_LOGIC;
		    BOT_Q: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE ALGO OF ffdh IS
BEGIN

	    PROCESS (CLK)
			BEGIN
				IF RISING_EDGE (CLK) THEN
					IF HAB = '1' THEN
						BOT_Q <= D;
					END IF;
				END IF;
			END PROCESS;
			
END ALGO;
